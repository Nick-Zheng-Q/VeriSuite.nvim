typedef enum logic [1:0] { IDLE, RUN, DONE } state_t;

module test_enum;
  /*AUTOASCIIENUM*/
endmodule
